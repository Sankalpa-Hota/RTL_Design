module TB_D_FF;
   reg